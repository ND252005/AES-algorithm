/*
Đầu vào: 
- clk:
- reset:
- độ dài khóa
- độ dài từ
- 
- flag_in:
Đầu ra:
- 
- 
*/

`timescale 1ns/1ps

module KeyExpantion #(
    parameter KEY_LEN = 128,
    parameter NUMS_OF_ROUND = 10,
    parameter WORD_LEN = 32
) (
    input clk,
    input reset,
    input [KEY_LEN-1 : 0] Secret_key,
    input valid_in,
    output wire [(NUMS_OF_ROUND*KEY_LEN-1) : 0] key_expan,
    output wire [NUMS_OF_ROUND-1 : 0] valid_out
);
    wire [KEY_LEN-1:0] key_arr [0 : NUMS_OF_ROUND];
    wire [NUMS_OF_ROUND-1:0] subkey_valid_out;


//---Rcon table---
wire [WORD_LEN-1:0] Rcon [0:9];
assign Rcon[0] = 32'h01000000;
assign Rcon[1] = 32'h02000000;
assign Rcon[2] = 32'h04000000;
assign Rcon[3] = 32'h08000000;
assign Rcon[4] = 32'h10000000;
assign Rcon[5] = 32'h20000000;
assign Rcon[6] = 32'h40000000;
assign Rcon[7] = 32'h80000000;
assign Rcon[8] = 32'h1B000000;
assign Rcon[9] = 32'h36000000;

GenSubKey #(
    .KEY_LEN(KEY_LEN)
    ) FGSK (
    .clk(clk),
    .reset(reset),
    .Rcon(Rcon[0]),
    .data_in(Secret_key),
    .valid_in(valid_in),
    .data_out(key_arr[0]),
    .valid_out(subkey_valid_out[0])
);

genvar i;
generate
    for(i = 1; i < NUMS_OF_ROUND; i = i+1) begin : gen_subkeys
    wire [KEY_LEN-1:0] prev_subkey = key_arr[i-1];
    wire prev_valid = subkey_valid_out[i-1];
    GenSubKey #(
    .KEY_LEN(KEY_LEN)
    ) GSK_inst (
    .clk(clk),
    .reset(reset),
    .Rcon(Rcon[i]),
    .data_in(prev_subkey),
    .valid_in(prev_valid),
    .data_out(key_arr[i]),
    .valid_out(subkey_valid_out[i])
);
    end
endgenerate

assign key_expan = {
    key_arr[9],
    key_arr[8],
    key_arr[7],
    key_arr[6],
    key_arr[5],
    key_arr[4],
    key_arr[3],
    key_arr[2],
    key_arr[1],
    key_arr[0]
    };
assign valid_out = subkey_valid_out;
    
endmodule