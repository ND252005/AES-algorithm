/*
Đầu vào: 
- clk:
- reset:
- length: độ dài khóa
- data_in:
- flag_in:
Đầu ra:
- 
- 
*/

`timescale 1ns/1ns

module KeyExpantion (
    
);
    
endmodule