/*
Đầu vào: 
- clk:
- reset:
- độ dài khóa
- độ dài từ
- 
- flag_in:
Đầu ra:
- 
- 
*/

`timescale 1ns/1ps

module KeyExpantion #(
    parameter KEY_LEN = 128,
    parameter NUMS_OF_ROUND = 14,
    parameter WORD_LEN = 32
) (
    input clk,
    input reset,
    input [KEY_LEN-1 : 0] low_cipher_key,
    input valid_in,
    output wire [(NUMS_OF_ROUND*KEY_LEN-1) : 0] key_expan,
    output wire [NUMS_OF_ROUND-1 : 0] valid_out
);
    wire [KEY_LEN-1:0] key_arr [0 : NUMS_OF_ROUND];
    wire [NUMS_OF_ROUND-1:0] subkey_valid_out;


//---Rcon table---
wire [WORD_LEN-1:0] Rcon [0:9];
assign Rcon[0] = 32'h01000000;
assign Rcon[1] = 32'h02000000;
assign Rcon[2] = 32'h04000000;
assign Rcon[3] = 32'h08000000;
assign Rcon[4] = 32'h10000000;
assign Rcon[5] = 32'h20000000;
assign Rcon[6] = 32'h40000000;
// assign Rcon[7] = 32'h80000000;
// assign Rcon[8] = 32'h1B000000;
// assign Rcon[9] = 32'h36000000;

// Round 2
GenSubKey #(
    .KEY_LEN(KEY_LEN)
    ) GSK_round_2 (
    .clk(clk),
    .reset(reset),
    .opcode(0),
    .Rcon(Rcon[0]),
    .data_in(Secret_key),
    .valid_in(valid_in),
    .data_out(key_arr[0]),
    .valid_out(subkey_valid_out[0])
);

// Round 3
GenSubKey #(
    .KEY_LEN(KEY_LEN)
    ) GSK_round_3 (
    .clk(clk),
    .reset(reset),
    .opcode(1),
    .Rcon(Rcon[0]),
    .data_in(key_arr[0]),
    .valid_in(subkey_valid_out[0]),
    .data_out(key_arr[1]),
    .valid_out(subkey_valid_out[1])
);

// Round 4
GenSubKey #(
    .KEY_LEN(KEY_LEN)
    ) GSK_round_4 (
    .clk(clk),
    .reset(reset),
    .opcode(0),
    .Rcon(Rcon[1]),
    .data_in(key_arr[1]),
    .valid_in(subkey_valid_out[1]),
    .data_out(key_arr[2]),
    .valid_out(subkey_valid_out[2])
);

// Round 5
GenSubKey #(
    .KEY_LEN(KEY_LEN)
    ) GSK_round_5 (
    .clk(clk),
    .reset(reset),
    .opcode(1),
    .Rcon(Rcon[1]),
    .data_in(key_arr[2]),
    .valid_in(subkey_valid_out[2]),
    .data_out(key_arr[3]),
    .valid_out(subkey_valid_out[3])
);

// Round 6
GenSubKey #(
    .KEY_LEN(KEY_LEN)
    ) GSK_round_6 (
    .clk(clk),
    .reset(reset),
    .opcode(0),
    .Rcon(Rcon[2]),
    .data_in(key_arr[3]),
    .valid_in(subkey_valid_out[3]),
    .data_out(key_arr[4]),
    .valid_out(subkey_valid_out[4])
);

// Round 7
GenSubKey #(
    .KEY_LEN(KEY_LEN)
    ) GSK_round_7 (
    .clk(clk),
    .reset(reset),
    .opcode(1),
    .Rcon(Rcon[2]),
    .data_in(key_arr[4]),
    .valid_in(subkey_valid_out[4]),
    .data_out(key_arr[5]),
    .valid_out(subkey_valid_out[5])
);

// Round 8
GenSubKey #(
    .KEY_LEN(KEY_LEN)
    ) GSK_round_8 (
    .clk(clk),
    .reset(reset),
    .opcode(0),
    .Rcon(Rcon[3]),
    .data_in(key_arr[5]),
    .valid_in(subkey_valid_out[5]),
    .data_out(key_arr[6]),
    .valid_out(subkey_valid_out[6])
);

// Round 9
GenSubKey #(
    .KEY_LEN(KEY_LEN)
    ) GSK_round_9 (
    .clk(clk),
    .reset(reset),
    .opcode(1),
    .Rcon(Rcon[3]),
    .data_in(key_arr[6]),
    .valid_in(subkey_valid_out[6]),
    .data_out(key_arr[7]),
    .valid_out(subkey_valid_out[7])
);

// Round 10
GenSubKey #(
    .KEY_LEN(KEY_LEN)
    ) GSK_round_10 (
    .clk(clk),
    .reset(reset),
    .opcode(0),
    .Rcon(Rcon[4]),
    .data_in(key_arr[7]),
    .valid_in(subkey_valid_out[7]),
    .data_out(key_arr[8]),
    .valid_out(subkey_valid_out[8])
);

// Round 11
GenSubKey #(
    .KEY_LEN(KEY_LEN)
    ) GSK_round_11 (
    .clk(clk),
    .reset(reset),
    .opcode(1),
    .Rcon(Rcon[4]),
    .data_in(key_arr[8]),
    .valid_in(subkey_valid_out[8]),
    .data_out(key_arr[9]),
    .valid_out(subkey_valid_out[9])
);

// Round 12
GenSubKey #(
    .KEY_LEN(KEY_LEN)
    ) GSK_round_12 (
    .clk(clk),
    .reset(reset),
    .opcode(0),
    .Rcon(Rcon[5]),
    .data_in(key_arr[9]),
    .valid_in(subkey_valid_out[9]),
    .data_out(key_arr[10]),
    .valid_out(subkey_valid_out[10])
);

// Round 13
GenSubKey #(
    .KEY_LEN(KEY_LEN)
    ) GSK_round_13 (
    .clk(clk),
    .reset(reset),
    .opcode(1),
    .Rcon(Rcon[5]),
    .data_in(key_arr[10]),
    .valid_in(subkey_valid_out[10]),
    .data_out(key_arr[11]),
    .valid_out(subkey_valid_out[11])
);

// Round 14
GenSubKey #(
    .KEY_LEN(KEY_LEN)
    ) GSK_round_14 (
    .clk(clk),
    .reset(reset),
    .opcode(0),
    .Rcon(Rcon[6]),
    .data_in(key_arr[11]),
    .valid_in(subkey_valid_out[11]),
    .data_out(key_arr[12]),
    .valid_out(subkey_valid_out[12])
);


assign key_expan = {
    key_arr[12],
    key_arr[11],
    key_arr[10],
    key_arr[9],
    key_arr[8],
    key_arr[7],
    key_arr[6],
    key_arr[5],
    key_arr[4],
    key_arr[3],
    key_arr[2],
    key_arr[1],
    key_arr[0]
    };
assign valid_out = subkey_valid_out;
    
endmodule